LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY USING_IR IS
  GENERIC (
    RX_HIGH_COUNT_MAX: STD_LOGIC_VECTOR(11 DOWNTO 0) := X"FFF";
    RX_HIGH_COUNT_MIN: STD_LOGIC_VECTOR(11 DOWNTO 0) := X"190";
    RX_LOW_COUNT_MAX : STD_LOGIC_VECTOR(11 DOWNTO 0) := X"258";
    RX_THRESHOLD     : STD_LOGIC_VECTOR(11 DOWNTO 0) := X"640"
  );
  PORT (
    CLOCK_50 : IN  STD_LOGIC_VECTOR(0 DOWNTO 0);
    SW      : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
    LED     : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
    IRDA_RXD: IN  STD_LOGIC_VECTOR(0 DOWNTO 0);
    HEX0    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX1    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX2    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX3    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX4    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX5    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END USING_IR;

ARCHITECTURE MAIN OF USING_IR IS
  SIGNAL CLOCK_50M         : STD_LOGIC := '0';
  SIGNAL CLOCK_1M          : STD_LOGIC := '0';
  SIGNAL RX_IN             : STD_LOGIC := '0';
  TYPE RX_PHASE_TYPE IS (IDLE, RX);
  SIGNAL RX_PHASE_NEXT     : RX_PHASE_TYPE := IDLE;
  SIGNAL RX_PHASE          : RX_PHASE_TYPE := IDLE;
  SIGNAL RX_NODE           : STD_LOGIC_VECTOR( 1 DOWNTO 0) := (OTHERS => '0');
  SIGNAL RX_HIGH_COUNT_NEXT: STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0'); 
  SIGNAL RX_HIGH_COUNT     : STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0'); 
  SIGNAL RX_LOW_COUNT_NEXT : STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0'); 
  SIGNAL RX_LOW_COUNT      : STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0'); 
  SIGNAL RX_SAMPLING       : STD_LOGIC := '0';
  SIGNAL RX_FRAME_NEXT     : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
  SIGNAL RX_FRAME          : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
  SIGNAL RX_ERROR          : STD_LOGIC := '0';
  SIGNAL RX_DATA_CHECK     : STD_LOGIC := '0';
  SIGNAL RX_DATA_NEXT      : STD_LOGIC_VECTOR( 7 DOWNTO 0) := (OTHERS => '0');
  SIGNAL RX_DATA           : STD_LOGIC_VECTOR( 7 DOWNTO 0) := (OTHERS => '0');
  COMPONENT HEX_ENCODE IS
    PORT(
      I: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
      O: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
    );
  END COMPONENT;
  COMPONENT PLL IS
    PORT (
      REFCLK   : IN  STD_LOGIC := 'X'; -- CLK
      RST      : IN  STD_LOGIC := 'X'; -- RESET
      OUTCLK_0 : OUT STD_LOGIC         -- CLK
    );
  END COMPONENT;
BEGIN
  CLOCK_50M <= CLOCK_50(0);
  LED <= "0000000001" WHEN RX_PHASE = IDLE ELSE
         "0000000010" WHEN RX_PHASE = RX ELSE "1111111111";
  RX_IN <= IRDA_RXD(0);
  PLL_MAP: PLL PORT MAP (CLOCK_50M, '0', CLOCK_1M);
  ------------------------------------------------------------
  RX_PHASE_NEXT <= IDLE WHEN RX_ERROR = '1' ELSE
                   RX WHEN RX_PHASE = IDLE AND RX_NODE(0) = '0' ELSE RX_PHASE;
  RX_HIGH_COUNT_NEXT <= RX_HIGH_COUNT + '1' WHEN RX_PHASE = RX AND RX_NODE(1) = '1' ELSE (OTHERS => '0');
  RX_LOW_COUNT_NEXT <= RX_LOW_COUNT + '1' WHEN RX_PHASE = RX AND RX_NODE(1) = '0' ELSE (OTHERS => '0');
  RX_SAMPLING <= '1' WHEN RX_NODE(0) = '0' AND RX_NODE(1) = '1' AND RX_HIGH_COUNT > RX_HIGH_COUNT_MIN ELSE '0';
  RX_FRAME_NEXT <= RX_FRAME WHEN RX_SAMPLING = '0' ELSE
                   '1' & RX_FRAME(15 DOWNTO 1) WHEN RX_HIGH_COUNT > RX_THRESHOLD ELSE '0' & RX_FRAME(15 DOWNTO 1);
  RX_ERROR <= '1' WHEN RX_HIGH_COUNT = RX_HIGH_COUNT_MAX OR RX_LOW_COUNT = RX_LOW_COUNT_MAX ELSE '0';
  RX_DATA_CHECK <= '1' WHEN RX_HIGH_COUNT = RX_HIGH_COUNT_MAX AND (NOT RX_FRAME(15 DOWNTO 8)) = RX_FRAME(7 DOWNTO 0) ELSE '0';
  RX_DATA_NEXT <= RX_FRAME(7 DOWNTO 0) WHEN RX_DATA_CHECK = '1' ELSE RX_DATA;
  PROCESS(CLOCK_1M)
  BEGIN
    IF CLOCK_1M'EVENT AND CLOCK_1M = '1' THEN
      RX_NODE(0) <= RX_IN;
      RX_NODE(1) <= RX_NODE(0);
      RX_PHASE <= RX_PHASE_NEXT;   
      RX_HIGH_COUNT <= RX_HIGH_COUNT_NEXT;         
      RX_LOW_COUNT <= RX_LOW_COUNT_NEXT;         
      RX_FRAME <= RX_FRAME_NEXT;
      -- RX_SUCCESS <= RX_DATA_CHECK;
      RX_DATA <= RX_DATA_NEXT;
    END IF;
  END PROCESS;
  --------------------------------------------------------
  HEX_ENCODE_MAP0: HEX_ENCODE PORT MAP(RX_DATA(3 DOWNTO 0), HEX0);
  HEX_ENCODE_MAP1: HEX_ENCODE PORT MAP(RX_DATA(7 DOWNTO 4), HEX1);
  HEX_ENCODE_MAP2: HEX_ENCODE PORT MAP(RX_FRAME(3 DOWNTO 0), HEX2);
  HEX_ENCODE_MAP3: HEX_ENCODE PORT MAP(RX_FRAME(7 DOWNTO 4), HEX3);
  HEX_ENCODE_MAP4: HEX_ENCODE PORT MAP(RX_FRAME(11 DOWNTO 8), HEX4);
  HEX_ENCODE_MAP5: HEX_ENCODE PORT MAP(RX_FRAME(15 DOWNTO 12), HEX5);
END MAIN;
