LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY AND_1BIT IS 
  PORT (
    A: IN  STD_LOGIC_VECTOR(0 DOWNTO 0);
    B: IN  STD_LOGIC_VECTOR(0 DOWNTO 0);
    S: OUT STD_LOGIC_VECTOR(0 DOWNTO 0)
  );
END AND_1BIT;

ARCHITECTURE MAIN OF AND_1BIT IS
BEGIN
  S <= A AND B;
END MAIN;
