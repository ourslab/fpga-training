LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY USING_GPIO IS
  PORT (
    SW    : IN    STD_LOGIC_VECTOR( 9 DOWNTO 0);
    HEX0  : OUT   STD_LOGIC_VECTOR( 6 DOWNTO 0);
    HEX1  : OUT   STD_LOGIC_VECTOR( 6 DOWNTO 0);
    HEX2  : OUT   STD_LOGIC_VECTOR( 6 DOWNTO 0);
    HEX3  : OUT   STD_LOGIC_VECTOR( 6 DOWNTO 0);
    HEX4  : OUT   STD_LOGIC_VECTOR( 6 DOWNTO 0);
    HEX5  : OUT   STD_LOGIC_VECTOR( 6 DOWNTO 0);
    GPIO_0: INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    GPIO_1: INOUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END USING_GPIO;

ARCHITECTURE MAIN OF USING_GPIO IS
BEGIN
  HEX0 <= "1000000" WHEN GPIO_1(3 DOWNTO 0) = "0000" ELSE
          "1111001" WHEN GPIO_1(3 DOWNTO 0) = "0001" ELSE
          "0100100" WHEN GPIO_1(3 DOWNTO 0) = "0010" ELSE
          "0110000" WHEN GPIO_1(3 DOWNTO 0) = "0011" ELSE
          "0011001" WHEN GPIO_1(3 DOWNTO 0) = "0100" ELSE
          "0010010" WHEN GPIO_1(3 DOWNTO 0) = "0101" ELSE
          "0000010" WHEN GPIO_1(3 DOWNTO 0) = "0110" ELSE
          "1111000" WHEN GPIO_1(3 DOWNTO 0) = "0111" ELSE
          "0000000" WHEN GPIO_1(3 DOWNTO 0) = "1000" ELSE
          "0010000" WHEN GPIO_1(3 DOWNTO 0) = "1001" ELSE
          "0001000" WHEN GPIO_1(3 DOWNTO 0) = "1010" ELSE
          "0000011" WHEN GPIO_1(3 DOWNTO 0) = "1011" ELSE
          "1000110" WHEN GPIO_1(3 DOWNTO 0) = "1100" ELSE
          "0100001" WHEN GPIO_1(3 DOWNTO 0) = "1101" ELSE
          "0000110" WHEN GPIO_1(3 DOWNTO 0) = "1110" ELSE
          "0001110" WHEN GPIO_1(3 DOWNTO 0) = "1111" ELSE (OTHERS => '0');
  HEX1 <= "1000000" WHEN GPIO_1(7 DOWNTO 4) = "0000" ELSE
          "1111001" WHEN GPIO_1(7 DOWNTO 4) = "0001" ELSE
          "0100100" WHEN GPIO_1(7 DOWNTO 4) = "0010" ELSE
          "0110000" WHEN GPIO_1(7 DOWNTO 4) = "0011" ELSE
          "0011001" WHEN GPIO_1(7 DOWNTO 4) = "0100" ELSE
          "0010010" WHEN GPIO_1(7 DOWNTO 4) = "0101" ELSE
          "0000010" WHEN GPIO_1(7 DOWNTO 4) = "0110" ELSE
          "1111000" WHEN GPIO_1(7 DOWNTO 4) = "0111" ELSE
          "0000000" WHEN GPIO_1(7 DOWNTO 4) = "1000" ELSE
          "0010000" WHEN GPIO_1(7 DOWNTO 4) = "1001" ELSE
          "0001000" WHEN GPIO_1(7 DOWNTO 4) = "1010" ELSE
          "0000011" WHEN GPIO_1(7 DOWNTO 4) = "1011" ELSE
          "1000110" WHEN GPIO_1(7 DOWNTO 4) = "1100" ELSE
          "0100001" WHEN GPIO_1(7 DOWNTO 4) = "1101" ELSE
          "0000110" WHEN GPIO_1(7 DOWNTO 4) = "1110" ELSE
          "0001110" WHEN GPIO_1(7 DOWNTO 4) = "1111" ELSE (OTHERS => '0');
   GPIO_0(7 DOWNTO 0) <= SW(7 DOWNTO 0);
   GPIO_0(35 DOWNTO 8) <= (OTHERS => '0');
END MAIN;

